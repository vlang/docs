module main

struct Topic {
	title            string
	markdown_content string
	url              string
}

module main

struct Page {
	title   string
	content string
}

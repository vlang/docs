module main

struct Topic {
	title string
	url   string
}

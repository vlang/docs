module main

struct Topic {
	title            string
	markdown_content string
	id               string
	url              string
}
